module i3c_secondary_master #(
    parameter MAX_DEVICES = 8  // Maximum number of devices on the I3C bus
) (
    input  logic        clk,          // System clock
    input  logic        reset_n,      // Active-low reset
    inout  logic        sda,          // Serial Data Line
    output logic        scl,          // Serial Clock Line

    // Mastership Request Signals
    input  logic        request_mastership,  // Signal to request mastership
    output logic        master_granted,      // Signal indicating mastership granted

    // In-Band Interrupt (IBI) Signals
    input  logic        ibi_request,         // IBI request from a device
    output logic        ibi_ack,             // IBI acknowledgment

    // Slave Mode Address
    input  logic [6:0]  slave_address        // Assigned dynamic address
);

    // ----------------------------------------
    // Internal Signals
    // ----------------------------------------
    typedef enum logic [1:0] {
        SLAVE_MODE,
        MASTER_REQUEST,
        MASTER_MODE
    } state_t;

    state_t current_state, next_state;

    logic sda_out_en;        // Enable SDA driving
    logic sda_drive;         // Value to drive on SDA
    assign sda = sda_out_en ? sda_drive : 1'bz;

    logic scl_drive;         // Clock signal
    assign scl = scl_drive;

    typedef struct packed {
        logic [7:0] bcr;              // Bus Characteristics Register
        logic [7:0] dcr;              // Device Characteristics Register
        logic [7:0] lvr;              // Legacy Virtual Register
        logic [6:0] dynamic_address;  // Dynamic address assigned by master
    } device_info_t;

    device_info_t devices[MAX_DEVICES];  // Device information array
    int device_count;                    // Number of devices on the bus
    logic [7:0] temp_data;               // Temporary data for task use

    // ----------------------------------------
    // State Machine
    // ----------------------------------------
    always_ff @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            current_state <= SLAVE_MODE;
        end else begin
            current_state <= next_state;
        end
    end

    always_comb begin
        case (current_state)
            SLAVE_MODE: begin
                if (request_mastership)
                    next_state = MASTER_REQUEST;
                else
                    next_state = SLAVE_MODE;
            end

            MASTER_REQUEST: begin
                if (master_granted)
                    next_state = MASTER_MODE;
                else
                    next_state = MASTER_REQUEST;
            end

            MASTER_MODE: begin
                if (!request_mastership)
                    next_state = SLAVE_MODE;
                else
                    next_state = MASTER_MODE;
            end

            default: next_state = SLAVE_MODE;
        endcase
    end

    // ----------------------------------------
    // Slave Mode Operation
    // ----------------------------------------
    always_ff @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            ibi_ack <= 1'b0;
        end else if (current_state == SLAVE_MODE) begin
            if (detect_ibi()) begin
                ibi_ack <= 1'b1;  // Acknowledge IBI
            end else begin
                ibi_ack <= 1'b0;
            end
        end
    end

    function logic detect_ibi();
        // Check for IBI on the bus (SDA held low during idle by another device)
        return (sda == 1'b0 && scl == 1'b1);
    endfunction

    // ----------------------------------------
    // Request Mastership
    // ----------------------------------------
    always_ff @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            master_granted <= 1'b0;
        end else if (current_state == MASTER_REQUEST) begin
            // Send mastership request and wait for grant
            send_ccc_command(8'h06);  // MR (Mastership Request)
            wait_ack();
            master_granted <= 1'b1;
        end else begin
            master_granted <= 1'b0;
        end
    end

    // ----------------------------------------
    // Master Mode Operation
    // ----------------------------------------
    always_ff @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            device_count <= 0;  // Reset device count
        end else if (current_state == MASTER_MODE) begin
            // Assign dynamic addresses and collect device info
            assign_dynamic_addresses();
            collect_device_info();
        end
    end

    // ----------------------------------------
    // Dynamic Address Assignment
    // ----------------------------------------
    task assign_dynamic_addresses();
        int i;
        automatic logic [6:0] dynamic_addr = 7'h10;
        for (i = 0; i < MAX_DEVICES; i++) begin
            receive_data(temp_data);
            devices[i].bcr = temp_data;

            receive_data(temp_data);
            devices[i].dcr = temp_data;

            receive_data(temp_data);
            devices[i].lvr = temp_data;

            devices[i].dynamic_address = dynamic_addr;
            dynamic_addr++;
        end
    endtask

    // ----------------------------------------
    // Collect Device Information
    // ----------------------------------------
    task collect_device_info();
        int i;
        for (i = 0; i < device_count; i++) begin
            receive_data(temp_data);
            devices[i].bcr = temp_data;

            receive_data(temp_data);
            devices[i].dcr = temp_data;

            receive_data(temp_data);
            devices[i].lvr = temp_data;
        end
    endtask

    // ----------------------------------------
    // Data Transfer Tasks
    // ----------------------------------------
    task send_ccc_command(input logic [7:0] ccc_command);
        // Send a Common Command Code (CCC)
        send_data(ccc_command);
    endtask

    task send_data(input logic [7:0] data);
        integer i;
        for (i = 7; i >= 0; i--) begin
            sda_drive <= data[i];
            sda_out_en <= 1'b1;
            @(posedge scl);
        end
        sda_out_en <= 1'b0;
    endtask

    task receive_data(output logic [7:0] data);
        integer i;
        for (i = 7; i >= 0; i--) begin
            @(posedge scl);
            data[i] = sda;
        end
    endtask

    task wait_ack();
        @(negedge scl);
        if (sda != 1'b0) $fatal("ACK not received!");
    endtask

endmodule
